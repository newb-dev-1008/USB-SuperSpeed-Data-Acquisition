----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Tue Apr 26 12:17:20 2022
-- Parameters for COREAHBTOAPB3
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 16;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant testbench : string( 1 to 4 ) := "User";
end coreparameters;
