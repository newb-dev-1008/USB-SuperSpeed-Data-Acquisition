-- D Flip Flop with Asynchronous Reset and Clock Enable
